module sim_emac;
tb_emac tb();
`include "tc_miim.v"
endmodule
