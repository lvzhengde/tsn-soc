module sim_emac;
tb_emac tb();
`include "tc_full_duplex_receive_1000M.v"
endmodule
